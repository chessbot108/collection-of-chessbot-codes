b0VIM 8.2      P�^�J ��  weiming                                 weiming-Q505UAR                         ~weiming/collection-of-chessbot-codes/codes/HDU/HDU_4614.cpp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 utf-8 3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           �                            U       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ad  B   �     �       �  �  �  �  �  �    j  X  F  7  (      �  �  �  �  �  �  �  p  U  ?  )      �  �  �  �  r  q  L    �  �  �  �  �  �  |  l  \  P  9  6    �  �  �  l    �
  �
  �
  a
  [
  W
  T
  >
  
  
  
  �	  �	  r	  V	  >	  
	  �  �  �  �  �  �  �  c  T  P  M    �  �  �  n  S        �  �  |  e  V  P  8    �  �  �  �  �  �  �  �  �  ^  3    �  �  �  �  e  $    �  �  �  �  �  �  �  �  y  P  J  E      �  �  �  �  �  �  �                                                                          for(int i = 0; i<(this->n - 1) + this->s; i++){     void print(){      }       return dq;       G(l, r, 0, 0, this->n, dq);       deque<int> dq;     deque<int> get_intervals(int l, int r){          }       return Q_sum(l, r, 0, 0, this->n);     long long query_sum(int l, int r){      }       S(l, r, 0, val, 0, this->n);     void set_val(int l, int r, int val){       }       }         siz[i] = siz[LC(i)] * 2;         arr[i] = make_pair(arr[LC(i)].first, arr[RC(i)].second);       for(int i = n - 2; i >= 0; i--){       }         siz[i] = 1;         arr[i] = make_pair(i - (n - 1), i - (n - 2));       for(int i = n - 1; i < n*2; i++){       memset(marked, false, sizeof(marked));       memset(set_tag, 0, sizeof(set_tag));       memset(sum, 0, sizeof(sum));       this->n = pow_2(LOG2(s));       this->s = s;     seg_tree(int s){    public:    }     G(qL, qR, RC(k), mid, R, dq);     G(qL, qR, LC(k), L, mid, dq);     int mid = (L + R) / 2;     push_down(k, L, R);     }       return ;       dq.push_back(k);     if(qL <= L && R <= qR){     if(R <= L || R <= qL || qR <= L) return;   void G(int qL, int qR, int k, int L, int R, deque<int>& dq){      }     return Q_sum(qL, qR, LC(k), L, mid) + Q_sum(qL, qR, RC(k), mid, R);     int mid = (L + R) / 2;     push_down(k, L, R);     if(qL <= L && R <= qR) return sum[k];     if(R <= L || R <= qL || qR <= L) return 0LL;     //printf("%d %d %d %d %d\n", qL, qR, k, L, R);   long long Q_sum(int qL, int qR, int k, int L, int R){       }     update(k);     S(qL, qR, RC(k), val, mid, R);     S(qL, qR, LC(k), val, L, mid);     int mid = (L + R) / 2;     push_down(k, L, R);      }       return ;       marked[k] = true;       sum[k] = (long long)val * (long long)(R - L);       set_tag[k] = val;     if(qL <= L && R <= qR){     if(R <= L || R <= qL || qR <= L) return;      //printf("%d %d %d %d %d %d\n", qL, qR, k, val, L, R);   void S(int qL, int qR, int k, int val, int L, int R){    }     sum[k] = sum[LC(k)] + sum[RC(k)];   void update(int k){      }     }       marked[LC(k)] = marked[RC(k)] = true; //mark       marked[k] = false; //reset mark       set_tag[k] = 0; //reset tag       sum[RC(k)] = (long long)(R - mid) * (long long)set_tag[k];        sum[LC(k)] = (long long)(mid - L) * (long long)set_tag[k]; //merge sums       int mid = (L + R) / 2;        set_tag[LC(k)] = set_tag[RC(k)] = set_tag[k]; //merge tag     if(marked[k]){     if(L + 1 == R) return; //nothing to push down   void push_down(int k, int L, int R){      //d is min, t is max   int s, n; class seg_tree{ int siz[max_v]; pair<int, int> arr[220000];   bool marked[max_v]; long long sum[max_v]; int set_tag[max_v], add[max_v];  } 	freopen((file_name+".out").c_str(), "w+", stdout); 	freopen((file_name+".in").c_str(), "r", stdin); void setIO(const string& file_name){  using namespace std; #define LOG2(n) ((int)ceil(log2((n)))) #define RC(n) (((n) << 1) + 2) #define LC(n) (((n) << 1) + 1) #define lsb(n) ((n)&(-(n))) //tree #define pow_2(n) (1 << n) #define byte_max 0x3f #define cont continue #define int_max 0x3f3f3f3f #define max_v 410000  #include <functional> //#include <unordered_set> //#include <unordered_map> #include <deque> #include <stack> #include <queue> #include <list> #include <sstream> #include <set> #include <map> #include <string> #include <vector> #include <algorithm> #include <cassert> #include <cmath> #include <ctime> #include <cstdlib> #include <cstring> #include <cstdio> #include <iostream> ad  �  	     U       T  L  <  6  1  .  -    �  �  �  r  C     �  �  �  �  �  �  ~  h  @    �  �  �  �  �  �  Y  J  4    �  �  J  �
  �
  �
  �
  �
  �
  �
  �
  �
  |
  n
  `
  E
  2
  
  	
  �	  �	  �	  �	  �	  o	  S	  	  �  �  �  {  D  6    �  �  �  �  �  �  �  T  8  0  *          
  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              } 	return 0;    }     puts("");     }       }         S.set_val(a, b, 0);         printf("O:%lld\n", S.query_sum(a, b));         b++;       }else{          }           S.set_val(L, R, 1);           printf("O:%d %d\n", L, R);           assert(R >= 0);           //if(R < 0) R = right_0(temp, R * -1);         else{         if(L == -1) printf("Can not take any one.\n");        // assert((L != -1) ^ (R != -1));         int R = right_0(temp, b);// puts("");         int L = left_0(temp);// puts("");        // puts("");        //   printf("%d, %d %d\n", X, arr[X].first, arr[X].second);        // for(int X : temp)         deque<int> temp = S.get_intervals(a, n);       if(t == 1){       S.print();       scanf("%d%d%d", &t, &a, &b);       int t, a, b;     while(q--){    // S.print();     S.set_val(0, n, 0);     seg_tree S(n);     scanf("%d%d", &n, &q);     int n, q;   while(T--){   scanf("%d", &T);   int T; int main(){   }   return DIE(DQ);   }     else dq.push_front(RC(cur)), dq.push_front(LC(cur));     else if(tot + 1 == b && sum[cur] == 0 && siz[cur] == 1) return arr[cur].first;     if(tot + siz[cur] - (int)sum[cur] < b) tot += siz[cur] -(int)sum[cur];  //   printf("%d, %d %d %d %lld\n", cur, arr[cur].first, arr[cur].second, siz[cur], sum[cur]);     int cur = dq.front(); dq.pop_front();   while(!dq.empty()){   deque<int> dq = DQ;   int tot = 0; int right_0(const deque<int>& DQ, int b){  }   return -1;   }     else dq.push_back(LC(cur)), dq.push_back(RC(cur));     else if(siz[cur] == 1 && sum[cur] == 0) return arr[cur].first;     if(marked[cur] && set_tag[cur] == 1) cont;     int cur = dq.back(); dq.pop_back();   while(!dq.empty()){   deque<int> dq = DQ; int DIE(const deque<int>& DQ){  }   return -1;   }     else dq.push_front(RC(cur)), dq.push_front(LC(cur));     else if(siz[cur] == 1 && sum[cur] == 0) return arr[cur].first;     if(marked[cur] && set_tag[cur] == 1) cont; //    printf("%d, %d %d\n", cur, arr[cur].first, arr[cur].second);     int cur = dq.front(); dq.pop_front();   while(!dq.empty()){   deque<int> dq = DQ; int left_0(const deque<int>& DQ){  };          }       puts("");       }         printf("%d:\n\tlc->%d, rc->%d\n\tleft_bound->%d, right_bound->%d\n\tsum->%lld\n\tset_tag->%d\n", i, LC(i), RC(i), arr[i].first, arr[i].second, sum[i], set_tag[i]); 